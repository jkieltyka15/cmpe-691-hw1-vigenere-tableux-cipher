module vtc_tb();

initial
  begin
    $display("Hello World!");
    $finish;
  end

endmodule